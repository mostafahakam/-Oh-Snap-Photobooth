// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7−0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDG7−0 are parallel port outputs from the Nios II system
module lights (SW, KEY, CLOCK_50, LEDR, DRAM_CLK, DRAM_CKE,
DRAM_ADDR, DRAM_BA, DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N,
DRAM_WE_N, DRAM_DQ, DRAM_UDQM, DRAM_LDQM, GPIO_0, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5);
input [7:0] SW;
input [2:0] KEY;
input CLOCK_50;
output [7:0] LEDR;
output [11:0] DRAM_ADDR;
output [1:0] DRAM_BA;
output DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK;
output DRAM_CKE, DRAM_CS_N, DRAM_WE_N, DRAM_UDQM, DRAM_LDQM;
inout [15:0] DRAM_DQ;
inout [35:0] GPIO_0;
output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;

wire RS232_rxd;
wire RS232_txd;
wire[19:0] sev_seg_export;

assign RS232_rxd = GPIO_0[34]; 
assign GPIO_0[32] = RS232_txd;

wire[3:0] hex_export0, hex_export1, hex_export2, hex_export3, hex_export4, hex_export5;

sev s0(hex_export0, HEX0);
sev s1(hex_export1, HEX1);
sev s2(hex_export2, HEX2);
sev s3(hex_export3, HEX3);
sev s4(hex_export4, HEX4);
sev s5(hex_export5, HEX5);


// Instantiate the Nios II system module generated by the Qsys tool:

tut_nios NoisII (
		.clk_clk(CLOCK_50),        //      clk_1.clk
		.leds_export(LEDR),      //       leds.export
		.reset_reset(~KEY[0]),    //    reset_1.reset
		.sdram_clk_clk(DRAM_CLK),    //  sdram_clk.clk
		.sdram_wire_addr(DRAM_ADDR),  // sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),    //           .ba
		.sdram_wire_cas_n(DRAM_CAS_N), //           .cas_n
		.sdram_wire_cke(DRAM_CKE),   //           .cke
		.sdram_wire_cs_n(DRAM_CS_N),  //           .cs_n
		.sdram_wire_dq(DRAM_DQ),    //           .dq
		.sdram_wire_dqm({DRAM_UDQM, DRAM_LDQM}),   //           .dqm
		.sdram_wire_ras_n(DRAM_RAS_N), //           .ras_n
		.sdram_wire_we_n(DRAM_WE_N),  //           .we_n
		.switches_export(SW),   //   switches.export
		.uart_rxd(RS232_rxd),         //       uart.rxd
		.uart_txd(RS232_txd),
		.pushbutton_export(~KEY[1]),
		.hex0_export(hex_export0),       //       hex0.export
		.hex1_export(hex_export1),       //       hex1.export
		.hex2_export(hex_export2),       //       hex2.export
		.hex3_export(hex_export3),       //       hex3.export
		.hex4_export(hex_export4),       //       hex4.export
		.hex5_export(hex_export5),       //       hex5.export		
	);
	

endmodule
