// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7−0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDG7−0 are parallel port outputs from the Nios II system
module lights (SW, KEY, CLOCK_50, LEDR, DRAM_CLK, DRAM_CKE,
DRAM_ADDR, DRAM_BA, DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N,
DRAM_WE_N, DRAM_DQ, DRAM_UDQM, DRAM_LDQM);
input [7:0] SW;
input [0:0] KEY;
input CLOCK_50;
output [7:0] LEDR;
output [11:0] DRAM_ADDR;
output [1:0] DRAM_BA;
output DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK;
output DRAM_CKE, DRAM_CS_N, DRAM_WE_N, DRAM_UDQM, DRAM_LDQM;
inout [15:0] DRAM_DQ;
// Instantiate the Nios II system module generated by the Qsys tool:

tut_nios NoisII (
		.clk_clk(CLOCK_50),        //      clk_1.clk
		.leds_export(LEDR),      //       leds.export
		.reset_reset(~KEY),    //    reset_1.reset
		.sdram_clk_clk(DRAM_CLK),    //  sdram_clk.clk
		.sdram_wire_addr(DRAM_ADDR),  // sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),    //           .ba
		.sdram_wire_cas_n(DRAM_CAS_N), //           .cas_n
		.sdram_wire_cke(DRAM_CKE),   //           .cke
		.sdram_wire_cs_n(DRAM_CS_N),  //           .cs_n
		.sdram_wire_dq(DRAM_DQ),    //           .dq
		.sdram_wire_dqm({DRAM_UDQM, DRAM_LDQM}),   //           .dqm
		.sdram_wire_ras_n(DRAM_RAS_N), //           .ras_n
		.sdram_wire_we_n(DRAM_WE_N),  //           .we_n
		.switches_export(SW)   //   switches.export
	);
	

endmodule
